//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: io_bottom]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Aug  8 10:08:34 2022
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

// ----- BEGIN Grid Verilog module: grid_io_bottom_bottom -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for grid_io_bottom_bottom -----
module grid_io_bottom_bottom(IO_ISOL_N,
                             config_readback,
                             config_enable,
                             pReset,
                             prog_clk,
                             gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN,
                             gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT,
                             gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR,
                             top_width_0_height_0_subtile_0__pin_outpad_0_,
                             top_width_0_height_0_subtile_1__pin_outpad_0_,
                             top_width_0_height_0_subtile_2__pin_outpad_0_,
                             top_width_0_height_0_subtile_3__pin_outpad_0_,
                             top_width_0_height_0_subtile_4__pin_outpad_0_,
                             top_width_0_height_0_subtile_5__pin_outpad_0_,
                             top_width_0_height_0_subtile_6__pin_outpad_0_,
                             top_width_0_height_0_subtile_7__pin_outpad_0_,
                             top_width_0_height_0_subtile_8__pin_outpad_0_,
                             ccff_head,
                             top_width_0_height_0_subtile_0__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_0__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_1__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_1__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_2__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_2__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_3__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_3__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_4__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_4__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_5__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_5__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_6__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_6__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_7__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_7__pin_inpad_0_lower,
                             top_width_0_height_0_subtile_8__pin_inpad_0_upper,
                             top_width_0_height_0_subtile_8__pin_inpad_0_lower,
                             ccff_tail);
//----- GLOBAL PORTS -----
input wire [0:0] IO_ISOL_N;
//----- GLOBAL PORTS -----
input wire [0:0] config_readback;
//----- GLOBAL PORTS -----
input wire [0:0] config_enable;
//----- GLOBAL PORTS -----
input wire [0:0] pReset;
//----- GLOBAL PORTS -----
input wire [0:0] prog_clk;
//----- GPIN PORTS -----
input wire [0:8] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN;
//----- GPOUT PORTS -----
output wire [0:8] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT;
//----- GPOUT PORTS -----
output wire [0:8] gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_0__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_1__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_2__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_3__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_4__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_5__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_6__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_7__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] top_width_0_height_0_subtile_8__pin_outpad_0_;
//----- INPUT PORTS -----
input wire [0:0] ccff_head;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_0__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_0__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_1__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_1__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_2__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_2__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_3__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_3__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_4__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_4__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_5__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_5__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_6__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_6__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_7__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_7__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_8__pin_inpad_0_upper;
//----- OUTPUT PORTS -----
output wire [0:0] top_width_0_height_0_subtile_8__pin_inpad_0_lower;
//----- OUTPUT PORTS -----
output wire [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] logical_tile_io_mode_io__0_ccff_tail;
wire [0:0] logical_tile_io_mode_io__1_ccff_tail;
wire [0:0] logical_tile_io_mode_io__2_ccff_tail;
wire [0:0] logical_tile_io_mode_io__3_ccff_tail;
wire [0:0] logical_tile_io_mode_io__4_ccff_tail;
wire [0:0] logical_tile_io_mode_io__5_ccff_tail;
wire [0:0] logical_tile_io_mode_io__6_ccff_tail;
wire [0:0] logical_tile_io_mode_io__7_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
	assign top_width_0_height_0_subtile_0__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_0__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_1__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_1__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_2__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_2__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_3__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_3__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_4__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_4__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_5__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_5__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_6__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_6__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_7__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_7__pin_inpad_0_upper[0];
	assign top_width_0_height_0_subtile_8__pin_inpad_0_lower[0] = top_width_0_height_0_subtile_8__pin_inpad_0_upper[0];
// ----- END Local output short connections -----

	logical_tile_io_mode_io_ logical_tile_io_mode_io__0 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[0]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[0]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[0]),
		.io_outpad(top_width_0_height_0_subtile_0__pin_outpad_0_),
		.ccff_head(ccff_head),
		.io_inpad(top_width_0_height_0_subtile_0__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__0_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__1 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[1]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[1]),
		.io_outpad(top_width_0_height_0_subtile_1__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__0_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_1__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__1_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__2 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[2]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[2]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[2]),
		.io_outpad(top_width_0_height_0_subtile_2__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__1_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_2__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__2_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__3 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[3]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[3]),
		.io_outpad(top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__2_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_3__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__3_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__4 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[4]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[4]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[4]),
		.io_outpad(top_width_0_height_0_subtile_4__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__3_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_4__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__4_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__5 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[5]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[5]),
		.io_outpad(top_width_0_height_0_subtile_5__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__4_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_5__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__5_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__6 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[6]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[6]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[6]),
		.io_outpad(top_width_0_height_0_subtile_6__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__5_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_6__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__6_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__7 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[7]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[7]),
		.io_outpad(top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__6_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_7__pin_inpad_0_upper),
		.ccff_tail(logical_tile_io_mode_io__7_ccff_tail));

	logical_tile_io_mode_io_ logical_tile_io_mode_io__8 (
		.IO_ISOL_N(IO_ISOL_N),
		.config_readback(config_readback),
		.config_enable(config_enable),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_IN[8]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_OUT[8]),
		.gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR(gfpga_pad_EMBEDDED_IO_ISOLN_SOC_DIR[8]),
		.io_outpad(top_width_0_height_0_subtile_8__pin_outpad_0_),
		.ccff_head(logical_tile_io_mode_io__7_ccff_tail),
		.io_inpad(top_width_0_height_0_subtile_8__pin_inpad_0_upper),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_io_bottom_bottom -----

//----- Default net type -----
`default_nettype none



// ----- END Grid Verilog module: grid_io_bottom_bottom -----

