

module pmu_top;




endmodule
